// megafunction wizard: %RAM: 2-PORT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altsyncram 

// ============================================================
// File Name: ram_dp_533.v
// Megafunction Name(s):
// 			altsyncram
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 11.1 Build 259 01/25/2012 SP 2 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module ram_dp_533 (
	address_a,
	address_b,
	clock,
	data_a,
	data_b,
	wren_a,
	wren_b,
	q_a,
	q_b);

	input	[17:0]  address_a;
	input	[17:0]  address_b;
	input	  clock;
	input	[7:0]  data_a;
	input	[7:0]  data_b;
	input	  wren_a;
	input	  wren_b;
	output	[7:0]  q_a;
	output	[7:0]  q_b;
//`ifndef ALTERA_RESERVED_QIS
//// synopsys translate_off
//`endif
//	tri1	  clock;
//	tri0	  wren_a;
//	tri0	  wren_b;
//`ifndef ALTERA_RESERVED_QIS
//// synopsys translate_on
//`endif

	wire [7:0] sub_wire0;
	wire [7:0] sub_wire1;
	wire [7:0] q_a = data_a[7:0];
	wire [7:0] q_b = sub_wire1[7:0];



//ram2 inst_ram2 (
//  .clka(clock),    // input wire clka
//  .wea(wren_a),      // input wire [0 : 0] wea
//  .addra(address_a),  // input wire [17 : 0] addra
//  .dina(data_a),    // input wire [7 : 0] dina
//  .douta(sub_wire0),  // output wire [7 : 0] douta
//  
//  .clkb(clock),    // input wire clkb
//  .web(wren_b),      // input wire [0 : 0] web
//  .addrb(address_b),  // input wire [17 : 0] addrb
//  .dinb(data_b),    // input wire [7 : 0] dinb
//  .doutb(sub_wire1)  // output wire [7 : 0] doutb
//);

ram2 inst_ram2 (
  .clka(clock),    // input wire clka
  .wea(wren_a),      // input wire [0 : 0] wea
  .addra(address_a),  // input wire [17 : 0] addra
  .dina(data_a),    // input wire [7 : 0] dina
  
  .clkb(clock),    // input wire clkb
  .enb(1'b1),      // input wire enb
  .addrb(address_b),  // input wire [17 : 0] addrb
  .doutb(sub_wire1)  // output wire [7 : 0] doutb
);




	//altsyncram	altsyncram_component (
	//			.clock0 (clock),
	//			.wren_a (wren_a),
	//			.address_b (address_b),
	//			.data_b (data_b),
	//			.wren_b (wren_b),
	//			.address_a (address_a),
	//			.data_a (data_a),
	//			.q_a (sub_wire0),
	//			.q_b (sub_wire1),
	//			.aclr0 (1'b0),
	//			.aclr1 (1'b0),
	//			.addressstall_a (1'b0),
	//			.addressstall_b (1'b0),
	//			.byteena_a (1'b1),
	//			.byteena_b (1'b1),
	//			.clock1 (1'b1),
	//			.clocken0 (1'b1),
	//			.clocken1 (1'b1),
	//			.clocken2 (1'b1),
	//			.clocken3 (1'b1),
	//			.eccstatus (),
	//			.rden_a (1'b1),
	//			.rden_b (1'b1));
	//defparam
	//	altsyncram_component.address_reg_b = "CLOCK0",
	//	altsyncram_component.clock_enable_input_a = "BYPASS",
	//	altsyncram_component.clock_enable_input_b = "BYPASS",
	//	altsyncram_component.clock_enable_output_a = "BYPASS",
	//	altsyncram_component.clock_enable_output_b = "BYPASS",
	//	altsyncram_component.indata_reg_b = "CLOCK0",
	//	altsyncram_component.intended_device_family = "Cyclone IV GX",
	//	altsyncram_component.lpm_type = "altsyncram",
	//	altsyncram_component.numwords_a = 213200,
	//	altsyncram_component.numwords_b = 213200,
	//	altsyncram_component.operation_mode = "BIDIR_DUAL_PORT",
	//	altsyncram_component.outdata_aclr_a = "NONE",
	//	altsyncram_component.outdata_aclr_b = "NONE",
	//	altsyncram_component.outdata_reg_a = "CLOCK0",
	//	altsyncram_component.outdata_reg_b = "CLOCK0",
	//	altsyncram_component.power_up_uninitialized = "FALSE",
	//	altsyncram_component.read_during_write_mode_mixed_ports = "DONT_CARE",
	//	altsyncram_component.read_during_write_mode_port_a = "NEW_DATA_NO_NBE_READ",
	//	altsyncram_component.read_during_write_mode_port_b = "NEW_DATA_NO_NBE_READ",
	//	altsyncram_component.widthad_a = 18,
	//	altsyncram_component.widthad_b = 18,
	//	altsyncram_component.width_a = 8,
	//	altsyncram_component.width_b = 8,
	//	altsyncram_component.width_byteena_a = 1,
	//	altsyncram_component.width_byteena_b = 1,
	//	altsyncram_component.wrcontrol_wraddress_reg_b = "CLOCK0";


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ADDRESSSTALL_A NUMERIC "0"
// Retrieval info: PRIVATE: ADDRESSSTALL_B NUMERIC "0"
// Retrieval info: PRIVATE: BYTEENA_ACLR_A NUMERIC "0"
// Retrieval info: PRIVATE: BYTEENA_ACLR_B NUMERIC "0"
// Retrieval info: PRIVATE: BYTE_ENABLE_A NUMERIC "0"
// Retrieval info: PRIVATE: BYTE_ENABLE_B NUMERIC "0"
// Retrieval info: PRIVATE: BYTE_SIZE NUMERIC "8"
// Retrieval info: PRIVATE: BlankMemory NUMERIC "1"
// Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_A NUMERIC "0"
// Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_B NUMERIC "0"
// Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_A NUMERIC "0"
// Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_B NUMERIC "0"
// Retrieval info: PRIVATE: CLRdata NUMERIC "0"
// Retrieval info: PRIVATE: CLRq NUMERIC "0"
// Retrieval info: PRIVATE: CLRrdaddress NUMERIC "0"
// Retrieval info: PRIVATE: CLRrren NUMERIC "0"
// Retrieval info: PRIVATE: CLRwraddress NUMERIC "0"
// Retrieval info: PRIVATE: CLRwren NUMERIC "0"
// Retrieval info: PRIVATE: Clock NUMERIC "0"
// Retrieval info: PRIVATE: Clock_A NUMERIC "0"
// Retrieval info: PRIVATE: Clock_B NUMERIC "0"
// Retrieval info: PRIVATE: ECC NUMERIC "0"
// Retrieval info: PRIVATE: ECC_PIPELINE_STAGE NUMERIC "0"
// Retrieval info: PRIVATE: IMPLEMENT_IN_LES NUMERIC "0"
// Retrieval info: PRIVATE: INDATA_ACLR_B NUMERIC "0"
// Retrieval info: PRIVATE: INDATA_REG_B NUMERIC "1"
// Retrieval info: PRIVATE: INIT_FILE_LAYOUT STRING "PORT_A"
// Retrieval info: PRIVATE: INIT_TO_SIM_X NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
// Retrieval info: PRIVATE: JTAG_ENABLED NUMERIC "0"
// Retrieval info: PRIVATE: JTAG_ID STRING "NONE"
// Retrieval info: PRIVATE: MAXIMUM_DEPTH NUMERIC "0"
// Retrieval info: PRIVATE: MEMSIZE NUMERIC "1705600"
// Retrieval info: PRIVATE: MEM_IN_BITS NUMERIC "0"
// Retrieval info: PRIVATE: MIFfilename STRING ""
// Retrieval info: PRIVATE: OPERATION_MODE NUMERIC "3"
// Retrieval info: PRIVATE: OUTDATA_ACLR_B NUMERIC "0"
// Retrieval info: PRIVATE: OUTDATA_REG_B NUMERIC "1"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
// Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_MIXED_PORTS NUMERIC "2"
// Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_A NUMERIC "3"
// Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_B NUMERIC "3"
// Retrieval info: PRIVATE: REGdata NUMERIC "1"
// Retrieval info: PRIVATE: REGq NUMERIC "1"
// Retrieval info: PRIVATE: REGrdaddress NUMERIC "0"
// Retrieval info: PRIVATE: REGrren NUMERIC "0"
// Retrieval info: PRIVATE: REGwraddress NUMERIC "1"
// Retrieval info: PRIVATE: REGwren NUMERIC "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: USE_DIFF_CLKEN NUMERIC "0"
// Retrieval info: PRIVATE: UseDPRAM NUMERIC "1"
// Retrieval info: PRIVATE: VarWidth NUMERIC "0"
// Retrieval info: PRIVATE: WIDTH_READ_A NUMERIC "8"
// Retrieval info: PRIVATE: WIDTH_READ_B NUMERIC "8"
// Retrieval info: PRIVATE: WIDTH_WRITE_A NUMERIC "8"
// Retrieval info: PRIVATE: WIDTH_WRITE_B NUMERIC "8"
// Retrieval info: PRIVATE: WRADDR_ACLR_B NUMERIC "0"
// Retrieval info: PRIVATE: WRADDR_REG_B NUMERIC "1"
// Retrieval info: PRIVATE: WRCTRL_ACLR_B NUMERIC "0"
// Retrieval info: PRIVATE: enable NUMERIC "0"
// Retrieval info: PRIVATE: rden NUMERIC "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: ADDRESS_REG_B STRING "CLOCK0"
// Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_A STRING "BYPASS"
// Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_B STRING "BYPASS"
// Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_A STRING "BYPASS"
// Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_B STRING "BYPASS"
// Retrieval info: CONSTANT: INDATA_REG_B STRING "CLOCK0"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altsyncram"
// Retrieval info: CONSTANT: NUMWORDS_A NUMERIC "213200"
// Retrieval info: CONSTANT: NUMWORDS_B NUMERIC "213200"
// Retrieval info: CONSTANT: OPERATION_MODE STRING "BIDIR_DUAL_PORT"
// Retrieval info: CONSTANT: OUTDATA_ACLR_A STRING "NONE"
// Retrieval info: CONSTANT: OUTDATA_ACLR_B STRING "NONE"
// Retrieval info: CONSTANT: OUTDATA_REG_A STRING "CLOCK0"
// Retrieval info: CONSTANT: OUTDATA_REG_B STRING "CLOCK0"
// Retrieval info: CONSTANT: POWER_UP_UNINITIALIZED STRING "FALSE"
// Retrieval info: CONSTANT: READ_DURING_WRITE_MODE_MIXED_PORTS STRING "DONT_CARE"
// Retrieval info: CONSTANT: READ_DURING_WRITE_MODE_PORT_A STRING "NEW_DATA_NO_NBE_READ"
// Retrieval info: CONSTANT: READ_DURING_WRITE_MODE_PORT_B STRING "NEW_DATA_NO_NBE_READ"
// Retrieval info: CONSTANT: WIDTHAD_A NUMERIC "18"
// Retrieval info: CONSTANT: WIDTHAD_B NUMERIC "18"
// Retrieval info: CONSTANT: WIDTH_A NUMERIC "8"
// Retrieval info: CONSTANT: WIDTH_B NUMERIC "8"
// Retrieval info: CONSTANT: WIDTH_BYTEENA_A NUMERIC "1"
// Retrieval info: CONSTANT: WIDTH_BYTEENA_B NUMERIC "1"
// Retrieval info: CONSTANT: WRCONTROL_WRADDRESS_REG_B STRING "CLOCK0"
// Retrieval info: USED_PORT: address_a 0 0 18 0 INPUT NODEFVAL "address_a[17..0]"
// Retrieval info: USED_PORT: address_b 0 0 18 0 INPUT NODEFVAL "address_b[17..0]"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT VCC "clock"
// Retrieval info: USED_PORT: data_a 0 0 8 0 INPUT NODEFVAL "data_a[7..0]"
// Retrieval info: USED_PORT: data_b 0 0 8 0 INPUT NODEFVAL "data_b[7..0]"
// Retrieval info: USED_PORT: q_a 0 0 8 0 OUTPUT NODEFVAL "q_a[7..0]"
// Retrieval info: USED_PORT: q_b 0 0 8 0 OUTPUT NODEFVAL "q_b[7..0]"
// Retrieval info: USED_PORT: wren_a 0 0 0 0 INPUT GND "wren_a"
// Retrieval info: USED_PORT: wren_b 0 0 0 0 INPUT GND "wren_b"
// Retrieval info: CONNECT: @address_a 0 0 18 0 address_a 0 0 18 0
// Retrieval info: CONNECT: @address_b 0 0 18 0 address_b 0 0 18 0
// Retrieval info: CONNECT: @clock0 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @data_a 0 0 8 0 data_a 0 0 8 0
// Retrieval info: CONNECT: @data_b 0 0 8 0 data_b 0 0 8 0
// Retrieval info: CONNECT: @wren_a 0 0 0 0 wren_a 0 0 0 0
// Retrieval info: CONNECT: @wren_b 0 0 0 0 wren_b 0 0 0 0
// Retrieval info: CONNECT: q_a 0 0 8 0 @q_a 0 0 8 0
// Retrieval info: CONNECT: q_b 0 0 8 0 @q_b 0 0 8 0
// Retrieval info: GEN_FILE: TYPE_NORMAL ram_dp_533.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram_dp_533.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram_dp_533.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram_dp_533.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram_dp_533_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram_dp_533_bb.v FALSE
// Retrieval info: LIB_FILE: altera_mf
