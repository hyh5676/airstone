// megafunction wizard: %LPM_MULT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altsquare 

// ============================================================
// File Name: mul5.v
// Megafunction Name(s):
// 			altsquare
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 11.1 Build 259 01/25/2012 SP 2 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module mul5 (
	aclr,
	clock,
	dataa,
	ena,
	result);

	input	  aclr;
	input	  clock;
	input	[20:0]  dataa;
	input	  ena;
	output	[41:0]  result;

	wire [41:0] sub_wire0;
	wire [41:0] result = sub_wire0[41:0];

	mult_5 inst_mult5 (
		.CLK(clock),    // input wire CLK
		.A(dataa),        // input wire [20 : 0] A
		.B(dataa),        // input wire [20 : 0] B
		.CE(ena),      // input wire CE
		.SCLR(aclr),  // input wire SCLR
		.P(sub_wire0)        // output wire [41 : 0] P
	);


	//altsquare	altsquare_component (
	//			.aclr (aclr),
	//			.clock (clock),
	//			.data (dataa),
	//			.ena (ena),
	//			.result (sub_wire0));
	//defparam
	//	altsquare_component.data_width = 21,
	//	altsquare_component.lpm_type = "ALTSQUARE",
	//	altsquare_component.pipeline = 2,
	//	altsquare_component.representation = "SIGNED",
	//	altsquare_component.result_width = 42;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: AutoSizeResult NUMERIC "1"
// Retrieval info: PRIVATE: B_isConstant NUMERIC "0"
// Retrieval info: PRIVATE: ConstantB NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix V"
// Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "2"
// Retrieval info: PRIVATE: Latency NUMERIC "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: SignedMult NUMERIC "1"
// Retrieval info: PRIVATE: USE_MULT NUMERIC "0"
// Retrieval info: PRIVATE: ValidConstant NUMERIC "0"
// Retrieval info: PRIVATE: WidthA NUMERIC "21"
// Retrieval info: PRIVATE: WidthB NUMERIC "8"
// Retrieval info: PRIVATE: WidthP NUMERIC "42"
// Retrieval info: PRIVATE: aclr NUMERIC "1"
// Retrieval info: PRIVATE: clken NUMERIC "1"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: PRIVATE: optimize NUMERIC "0"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: DATA_WIDTH NUMERIC "21"
// Retrieval info: CONSTANT: LPM_TYPE STRING "ALTSQUARE"
// Retrieval info: CONSTANT: PIPELINE NUMERIC "2"
// Retrieval info: CONSTANT: REPRESENTATION STRING "SIGNED"
// Retrieval info: CONSTANT: RESULT_WIDTH NUMERIC "42"
// Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL "aclr"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: dataa 0 0 21 0 INPUT NODEFVAL "dataa[20..0]"
// Retrieval info: USED_PORT: ena 0 0 0 0 INPUT NODEFVAL "ena"
// Retrieval info: USED_PORT: result 0 0 42 0 OUTPUT NODEFVAL "result[41..0]"
// Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 21 0 dataa 0 0 21 0
// Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
// Retrieval info: CONNECT: result 0 0 42 0 @result 0 0 42 0
// Retrieval info: GEN_FILE: TYPE_NORMAL mul.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL mul.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mul.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mul.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mul_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mul_bb.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL mul5.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL mul5.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mul5.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mul5.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mul5_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mul5_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
