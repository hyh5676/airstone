// megafunction wizard: %Shift register (RAM-based)%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSHIFT_TAPS 

// ============================================================
// File Name: line_buffer_31.v
// Megafunction Name(s):
// 			ALTSHIFT_TAPS
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 11.1 Build 259 01/25/2012 SP 2 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module line_buffer_31_571 (
	clken,
	clock,
	shiftin,
	shiftout,
	taps0x,
	taps10x,
	taps11x,
	taps12x,
	taps13x,
	taps14x,
	taps15x,
	taps16x,
	taps17x,
	taps18x,
	taps19x,
	taps1x,
	taps20x,
	taps21x,
	taps22x,
	taps23x,
	taps24x,
	taps25x,
	taps26x,
	taps27x,
	taps28x,
	taps29x,
	taps2x,
	taps30x,
	taps3x,
	taps4x,
	taps5x,
	taps6x,
	taps7x,
	taps8x,
	taps9x);

	input	  clken;
	input	  clock;
	input	[7:0]  shiftin;
	output	[7:0]  shiftout;
	output	[7:0]  taps0x ;
	output	[7:0]  taps10x;
	output	[7:0]  taps11x;
	output	[7:0]  taps12x;
	output	[7:0]  taps13x;
	output	[7:0]  taps14x;
	output	[7:0]  taps15x;
	output	[7:0]  taps16x;
	output	[7:0]  taps17x;
	output	[7:0]  taps18x;
	output	[7:0]  taps19x;
	output	[7:0]  taps1x ;
	output	[7:0]  taps20x;
	output	[7:0]  taps21x;
	output	[7:0]  taps22x;
	output	[7:0]  taps23x;
	output	[7:0]  taps24x;
	output	[7:0]  taps25x;
	output	[7:0]  taps26x;
	output	[7:0]  taps27x;
	output	[7:0]  taps28x;
	output	[7:0]  taps29x;
	output	[7:0]  taps2x ;
	output	[7:0]  taps30x;
	output	[7:0]  taps3x ;
	output	[7:0]  taps4x ;
	output	[7:0]  taps5x ;
	output	[7:0]  taps6x ;
	output	[7:0]  taps7x ;
	output	[7:0]  taps8x ;
	output	[7:0]  taps9x ;
	
	
	parameter tap_distance = 571;
    wire [7:0] taps_temp [0:31] ; // 32-bit array of wires
    reg  [31:0]clken_temp	; // 32-bit array of wires	
	reg [9:0]count;	

	wire [7:0] taps0x 	 =	 taps_temp[0 ];
	wire [7:0] taps10x   =   taps_temp[10];
	wire [7:0] taps11x   =   taps_temp[11];
	wire [7:0] taps12x   =   taps_temp[12];
	wire [7:0] taps13x   =   taps_temp[13];
	wire [7:0] taps14x   =   taps_temp[14];
	wire [7:0] taps15x   =   taps_temp[15];
	wire [7:0] taps16x   =   taps_temp[16];
	wire [7:0] taps17x   =   taps_temp[17];
	wire [7:0] taps18x   =   taps_temp[18];
	wire [7:0] taps19x   =   taps_temp[19];
	wire [7:0] taps1x   =   taps_temp[1 ];
	wire [7:0] taps20x   =   taps_temp[20];
	wire [7:0] taps21x   =   taps_temp[21];
	wire [7:0] taps22x   =   taps_temp[22];
	wire [7:0] taps23x   =   taps_temp[23];
	wire [7:0] taps24x   =   taps_temp[24];
	wire [7:0] taps25x   =   taps_temp[25];
	wire [7:0] taps26x   =   taps_temp[26];
	wire [7:0] taps27x   =   taps_temp[27];
	wire [7:0] taps28x   =   taps_temp[28];
	wire [7:0] taps29x   =   taps_temp[29];
	wire [7:0] taps2x   =   taps_temp[2 ];
	wire [7:0] taps30x   =   taps_temp[30];
	wire [7:0] taps3x   =   taps_temp[3 ];
	wire [7:0] taps4x   =   taps_temp[4 ];
	wire [7:0] taps5x   =   taps_temp[5 ];
	wire [7:0] taps6x   =   taps_temp[6 ];
	wire [7:0] taps7x   =   taps_temp[7 ];
	wire [7:0] taps8x   =   taps_temp[8 ];
	wire [7:0] taps9x   =   taps_temp[9 ];
	wire [7:0] shiftout  =   shiftin	  ;	



    always @(posedge clock) begin
		
        if (count == tap_distance-1 && clken) begin
            // Shift clk_temp array
            clken_temp[31:1] <= clken_temp[30:0]; // 将数组向左移位
            clken_temp[0] <= clken; // 将当前clk赋值到clk_temp[0]
			count <= 0;
        end
        else if(clken) begin
            count <= count + 1;
			clken_temp<=clken_temp;
		end
		else begin
            count <= 0;
			clken_temp<=0;		
		end
    end


    
    // Generate block for instantiating 32 instances of c_shift_ram_0
    genvar i;
    generate
        for (i = 0; i < 32; i = i + 1) begin : gen_inst_shift_ram
            c_shift_ram_0 inst_shift_ram (
                .A(tap_distance),    // input wire [9:0] A
                .D(i == 0 ? shiftin : taps_temp[i-1]), // input wire [7:0] D
                .CLK(clock),         // input wire CLK
                .CE(clken_temp[i]),          // input wire CE
                .Q(taps_temp[i])     // output wire [7:0] Q
            );
        end
    endgenerate


	//altshift_taps	ALTSHIFT_TAPS_component (
	//			.clock (clock),
	//			.clken (clken),
	//			.shiftin (shiftin),
	//			.taps (sub_wire0),
	//			.shiftout (sub_wire43),
	//			// synopsys translate_off,
	//			.aclr ()
	//			// synopsys translate_on
	//			);
	//defparam
	//	ALTSHIFT_TAPS_component.intended_device_family = "Cyclone IV GX",
	//	ALTSHIFT_TAPS_component.lpm_hint = "RAM_BLOCK_TYPE=AUTO",
	//	ALTSHIFT_TAPS_component.lpm_type = "altshift_taps",
	//	ALTSHIFT_TAPS_component.number_of_taps = 31,
	//	ALTSHIFT_TAPS_component.tap_distance = 678,
	//	ALTSHIFT_TAPS_component.width = 8;


endmodule

