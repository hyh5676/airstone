// megafunction wizard: %LPM_MULT%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_mult 

// ============================================================
// File Name: mul8.v
// Megafunction Name(s):
// 			lpm_mult
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 11.1 Build 259 01/25/2012 SP 2 SJ Full Version
// ************************************************************

//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module mul8 (
	aclr,
	clock,
	dataa,
	result);

	input	  aclr;
	input	  clock;
	input	[9:0]  dataa;
	output	[22:0]  result;

	wire [22:0] sub_wire0;	
	wire [12:0] sub_wire1 = 13'h1333;
	wire [22:0] result = sub_wire0[22:0];	
	
	mult_7 inst_mult8 (
		.CLK(clock),    // input wire CLK
		.A(dataa),        // input wire [9 : 0] A
		.B(sub_wire1),        // input wire [12 : 0] B
		.CE(1'b1),      // input wire CE
		.SCLR(aclr),  // input wire SCLR
		.P(sub_wire0)        // output wire [22 : 0] P
	);


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: AutoSizeResult NUMERIC "1"
// Retrieval info: PRIVATE: B_isConstant NUMERIC "1"
// Retrieval info: PRIVATE: ConstantB NUMERIC "4915"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix V"
// Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "5"
// Retrieval info: PRIVATE: Latency NUMERIC "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: SignedMult NUMERIC "0"
// Retrieval info: PRIVATE: USE_MULT NUMERIC "1"
// Retrieval info: PRIVATE: ValidConstant NUMERIC "1"
// Retrieval info: PRIVATE: WidthA NUMERIC "10"
// Retrieval info: PRIVATE: WidthB NUMERIC "13"
// Retrieval info: PRIVATE: WidthP NUMERIC "23"
// Retrieval info: PRIVATE: aclr NUMERIC "1"
// Retrieval info: PRIVATE: clken NUMERIC "0"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: PRIVATE: optimize NUMERIC "0"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_HINT STRING "INPUT_B_IS_CONSTANT=YES,MAXIMIZE_SPEED=5"
// Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "5"
// Retrieval info: CONSTANT: LPM_REPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MULT"
// Retrieval info: CONSTANT: LPM_WIDTHA NUMERIC "10"
// Retrieval info: CONSTANT: LPM_WIDTHB NUMERIC "13"
// Retrieval info: CONSTANT: LPM_WIDTHP NUMERIC "23"
// Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL "aclr"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: dataa 0 0 10 0 INPUT NODEFVAL "dataa[9..0]"
// Retrieval info: USED_PORT: result 0 0 23 0 OUTPUT NODEFVAL "result[22..0]"
// Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @dataa 0 0 10 0 dataa 0 0 10 0
// Retrieval info: CONNECT: @datab 0 0 13 0 4915 0 0 13 0
// Retrieval info: CONNECT: result 0 0 23 0 @result 0 0 23 0
// Retrieval info: GEN_FILE: TYPE_NORMAL mul8.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL mul8.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mul8.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mul8.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mul8_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mul8_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
