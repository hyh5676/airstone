// megafunction wizard: %ALTSQRT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSQRT 

// ============================================================
// File Name: sqrt.v
// Megafunction Name(s):
// 			ALTSQRT
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 11.1 Build 259 01/25/2012 SP 2 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module sqrt (
	aclr,
	clk,
	ena,
	radical,
	q,
	remainder);

	input	  aclr;
	input	  clk;
	input	  ena;
	input	[40:0]  radical;
	output	[20:0]  q;
	output	[21:0]  remainder;

	wire [20:0] sub_wire0;
	wire [0:0] sub_wire1;
	wire [20:0] q = sub_wire0[20:0];
	wire [21:0] remainder = sub_wire1;

	cordic_0 inst_cordic (
		.aclk(clk),                                        // input wire aclk
		.aclken(ena),                                    // input wire aclken
		.aresetn(~aclr),                                  // input wire aresetn
		.s_axis_cartesian_tvalid(ena),  // input wire s_axis_cartesian_tvalid
		.s_axis_cartesian_tdata(radical),    // input wire [47 : 0] s_axis_cartesian_tdata
		.m_axis_dout_tvalid(sub_wire1),            // output wire m_axis_dout_tvalid
		.m_axis_dout_tdata(sub_wire0)              // output wire [23 : 0] m_axis_dout_tdata
	);



	//altsqrt	ALTSQRT_component (
	//			.aclr (aclr),
	//			.clk (clk),
	//			.ena (ena),
	//			.radical (radical),
	//			.q (sub_wire0),
	//			.remainder (sub_wire1));
	//defparam
	//	ALTSQRT_component.pipeline = 16,
	//	ALTSQRT_component.q_port_width = 21,
	//	ALTSQRT_component.r_port_width = 22,
	//	ALTSQRT_component.width = 41;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: PIPELINE NUMERIC "16"
// Retrieval info: CONSTANT: Q_PORT_WIDTH NUMERIC "21"
// Retrieval info: CONSTANT: R_PORT_WIDTH NUMERIC "22"
// Retrieval info: CONSTANT: WIDTH NUMERIC "41"
// Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL "aclr"
// Retrieval info: USED_PORT: clk 0 0 0 0 INPUT NODEFVAL "clk"
// Retrieval info: USED_PORT: ena 0 0 0 0 INPUT NODEFVAL "ena"
// Retrieval info: USED_PORT: q 0 0 21 0 OUTPUT NODEFVAL "q[20..0]"
// Retrieval info: USED_PORT: radical 0 0 41 0 INPUT NODEFVAL "radical[40..0]"
// Retrieval info: USED_PORT: remainder 0 0 22 0 OUTPUT NODEFVAL "remainder[21..0]"
// Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
// Retrieval info: CONNECT: @clk 0 0 0 0 clk 0 0 0 0
// Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
// Retrieval info: CONNECT: @radical 0 0 41 0 radical 0 0 41 0
// Retrieval info: CONNECT: q 0 0 21 0 @q 0 0 21 0
// Retrieval info: CONNECT: remainder 0 0 22 0 @remainder 0 0 22 0
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
