// megafunction wizard: %Shift register (RAM-based)%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSHIFT_TAPS 

// ============================================================
// File Name: line_buffer_11_571.v
// Megafunction Name(s):
// 			ALTSHIFT_TAPS
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 11.1 Build 259 01/25/2012 SP 2 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module line_buffer_11_571 (
	clken,
	clock,
	shiftin,
	shiftout,
	taps0x,
	taps10x,
	taps1x,
	taps2x,
	taps3x,
	taps4x,
	taps5x,
	taps6x,
	taps7x,
	taps8x,
	taps9x);

	input	  clken;
	input	  clock;
	input	[7:0]  shiftin;
	output	[7:0]  shiftout;
	output	[7:0]  taps0x;
	output	[7:0]  taps10x;
	output	[7:0]  taps1x;
	output	[7:0]  taps2x;
	output	[7:0]  taps3x;
	output	[7:0]  taps4x;
	output	[7:0]  taps5x;
	output	[7:0]  taps6x;
	output	[7:0]  taps7x;
	output	[7:0]  taps8x;
	output	[7:0]  taps9x;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  clken;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire [87:0] sub_wire0;
	wire [7:0] sub_wire13;
	wire [63:56] sub_wire21 = sub_wire0[63:56];
	wire [31:24] sub_wire20 = sub_wire0[31:24];
	wire [31:24] sub_wire19 = sub_wire20[31:24];
	wire [55:48] sub_wire18 = sub_wire0[55:48];
	wire [55:48] sub_wire17 = sub_wire18[55:48];
	wire [23:16] sub_wire16 = sub_wire0[23:16];
	wire [23:16] sub_wire15 = sub_wire16[23:16];
	wire [79:72] sub_wire14 = sub_wire0[79:72];
	wire [79:72] sub_wire12 = sub_wire14[79:72];
	wire [47:40] sub_wire11 = sub_wire0[47:40];
	wire [47:40] sub_wire10 = sub_wire11[47:40];
	wire [15:8] sub_wire9 = sub_wire0[15:8];
	wire [15:8] sub_wire8 = sub_wire9[15:8];
	wire [87:80] sub_wire7 = sub_wire0[87:80];
	wire [87:80] sub_wire6 = sub_wire7[87:80];
	wire [71:64] sub_wire5 = sub_wire0[71:64];
	wire [71:64] sub_wire4 = sub_wire5[71:64];
	wire [39:32] sub_wire3 = sub_wire0[39:32];
	wire [39:32] sub_wire2 = sub_wire3[39:32];
	wire [7:0] sub_wire1 = sub_wire0[7:0];
	wire [7:0] taps0x = sub_wire1[7:0];
	wire [7:0] taps4x = sub_wire2[39:32];
	wire [7:0] taps8x = sub_wire4[71:64];
	wire [7:0] taps10x = sub_wire6[87:80];
	wire [7:0] taps1x = sub_wire8[15:8];
	wire [7:0] taps5x = sub_wire10[47:40];
	wire [7:0] taps9x = sub_wire12[79:72];
	wire [7:0] shiftout = sub_wire13[7:0];
	wire [7:0] taps2x = sub_wire15[23:16];
	wire [7:0] taps6x = sub_wire17[55:48];
	wire [7:0] taps3x = sub_wire19[31:24];
	wire [7:0] taps7x = sub_wire21[63:56];

	altshift_taps	ALTSHIFT_TAPS_component (
				.clock (clock),
				.clken (clken),
				.shiftin (shiftin),
				.taps (sub_wire0),
				.shiftout (sub_wire13)
				// synopsys translate_off
				,
				.aclr ()
				// synopsys translate_on
				);
	defparam
		ALTSHIFT_TAPS_component.intended_device_family = "Cyclone IV GX",
		ALTSHIFT_TAPS_component.lpm_hint = "RAM_BLOCK_TYPE=M9K",
		ALTSHIFT_TAPS_component.lpm_type = "altshift_taps",
		ALTSHIFT_TAPS_component.number_of_taps = 11,
		ALTSHIFT_TAPS_component.tap_distance = 571,
		ALTSHIFT_TAPS_component.width = 8;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACLR NUMERIC "0"
// Retrieval info: PRIVATE: CLKEN NUMERIC "1"
// Retrieval info: PRIVATE: GROUP_TAPS NUMERIC "1"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
// Retrieval info: PRIVATE: NUMBER_OF_TAPS NUMERIC "11"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: TAP_DISTANCE NUMERIC "571"
// Retrieval info: PRIVATE: WIDTH NUMERIC "8"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
// Retrieval info: CONSTANT: LPM_HINT STRING "RAM_BLOCK_TYPE=M9K"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altshift_taps"
// Retrieval info: CONSTANT: NUMBER_OF_TAPS NUMERIC "11"
// Retrieval info: CONSTANT: TAP_DISTANCE NUMERIC "571"
// Retrieval info: CONSTANT: WIDTH NUMERIC "8"
// Retrieval info: USED_PORT: clken 0 0 0 0 INPUT VCC "clken"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: shiftin 0 0 8 0 INPUT NODEFVAL "shiftin[7..0]"
// Retrieval info: USED_PORT: shiftout 0 0 8 0 OUTPUT NODEFVAL "shiftout[7..0]"
// Retrieval info: USED_PORT: taps0x 0 0 8 0 OUTPUT NODEFVAL "taps0x[7..0]"
// Retrieval info: USED_PORT: taps10x 0 0 8 0 OUTPUT NODEFVAL "taps10x[7..0]"
// Retrieval info: USED_PORT: taps1x 0 0 8 0 OUTPUT NODEFVAL "taps1x[7..0]"
// Retrieval info: USED_PORT: taps2x 0 0 8 0 OUTPUT NODEFVAL "taps2x[7..0]"
// Retrieval info: USED_PORT: taps3x 0 0 8 0 OUTPUT NODEFVAL "taps3x[7..0]"
// Retrieval info: USED_PORT: taps4x 0 0 8 0 OUTPUT NODEFVAL "taps4x[7..0]"
// Retrieval info: USED_PORT: taps5x 0 0 8 0 OUTPUT NODEFVAL "taps5x[7..0]"
// Retrieval info: USED_PORT: taps6x 0 0 8 0 OUTPUT NODEFVAL "taps6x[7..0]"
// Retrieval info: USED_PORT: taps7x 0 0 8 0 OUTPUT NODEFVAL "taps7x[7..0]"
// Retrieval info: USED_PORT: taps8x 0 0 8 0 OUTPUT NODEFVAL "taps8x[7..0]"
// Retrieval info: USED_PORT: taps9x 0 0 8 0 OUTPUT NODEFVAL "taps9x[7..0]"
// Retrieval info: CONNECT: @clken 0 0 0 0 clken 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @shiftin 0 0 8 0 shiftin 0 0 8 0
// Retrieval info: CONNECT: shiftout 0 0 8 0 @shiftout 0 0 8 0
// Retrieval info: CONNECT: taps0x 0 0 8 0 @taps 0 0 8 0
// Retrieval info: CONNECT: taps10x 0 0 8 0 @taps 0 0 8 80
// Retrieval info: CONNECT: taps1x 0 0 8 0 @taps 0 0 8 8
// Retrieval info: CONNECT: taps2x 0 0 8 0 @taps 0 0 8 16
// Retrieval info: CONNECT: taps3x 0 0 8 0 @taps 0 0 8 24
// Retrieval info: CONNECT: taps4x 0 0 8 0 @taps 0 0 8 32
// Retrieval info: CONNECT: taps5x 0 0 8 0 @taps 0 0 8 40
// Retrieval info: CONNECT: taps6x 0 0 8 0 @taps 0 0 8 48
// Retrieval info: CONNECT: taps7x 0 0 8 0 @taps 0 0 8 56
// Retrieval info: CONNECT: taps8x 0 0 8 0 @taps 0 0 8 64
// Retrieval info: CONNECT: taps9x 0 0 8 0 @taps 0 0 8 72
// Retrieval info: GEN_FILE: TYPE_NORMAL line_buffer_11_571.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL line_buffer_11_571.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL line_buffer_11_571.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL line_buffer_11_571.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL line_buffer_11_571_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL line_buffer_11_571_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
