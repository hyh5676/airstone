// megafunction wizard: %LPM_DIVIDE%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_DIVIDE 

// ============================================================
// File Name: div.v
// Megafunction Name(s):
// 			LPM_DIVIDE
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 11.1 Build 259 01/25/2012 SP 2 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module div (
	clock,
	denom,
	numer,
	quotient,
	remain);

	input	  clock;
	input	[20:0]  denom;
	input	[32:0]  numer;
	output	[32:0]  quotient;
	output	[20:0]  remain;

	//wire [20:0] sub_wire0;
	//wire [32:0] sub_wire1;
	wire [55 : 0] m_axis_dout_tdata;	
	wire [55 : 0] s_axis_divisor_tready,s_axis_dividend_tready;
	
	
	wire [20:0] remain = m_axis_dout_tdata[20:0];
	wire [32:0] quotient = m_axis_dout_tdata[53:21];


	div_gen_0 inst_div_gen (
		.aclk(clock),                                      // input wire aclk
		.aclken(1'b1),                                  // input wire aclken
		.aresetn(1'b1),                                // input wire aresetn
		.s_axis_divisor_tvalid(1'b1),    // input wire s_axis_divisor_tvalid
		.s_axis_divisor_tready(s_axis_divisor_tready),    // output wire s_axis_divisor_tready
		.s_axis_divisor_tdata(denom),      // input wire [23 : 0] s_axis_divisor_tdata
		.s_axis_dividend_tvalid(1'b1),  // input wire s_axis_dividend_tvalid
		.s_axis_dividend_tready(s_axis_dividend_tready),  // output wire s_axis_dividend_tready
		.s_axis_dividend_tdata(numer),    // input wire [39 : 0] s_axis_dividend_tdata
		.m_axis_dout_tvalid(m_axis_dout_tvalid),          // output wire m_axis_dout_tvalid
		.m_axis_dout_tdata(m_axis_dout_tdata)            // output wire [55 : 0] m_axis_dout_tdata
	);


	//lpm_divide	LPM_DIVIDE_component (
	//			.clock (clock),
	//			.denom (denom),
	//			.numer (numer),
	//			.remain (sub_wire0),
	//			.quotient (sub_wire1),
	//			.aclr (1'b0),
	//			.clken (1'b1));
	//defparam
	//	LPM_DIVIDE_component.lpm_drepresentation = "UNSIGNED",
	//	LPM_DIVIDE_component.lpm_hint = "LPM_REMAINDERPOSITIVE=TRUE",
	//	LPM_DIVIDE_component.lpm_nrepresentation = "SIGNED",
	//	LPM_DIVIDE_component.lpm_pipeline = 25,
	//	LPM_DIVIDE_component.lpm_type = "LPM_DIVIDE",
	//	LPM_DIVIDE_component.lpm_widthd = 21,
	//	LPM_DIVIDE_component.lpm_widthn = 33;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
// Retrieval info: PRIVATE: PRIVATE_LPM_REMAINDERPOSITIVE STRING "TRUE"
// Retrieval info: PRIVATE: PRIVATE_MAXIMIZE_SPEED NUMERIC "-1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: USING_PIPELINE NUMERIC "1"
// Retrieval info: PRIVATE: VERSION_NUMBER NUMERIC "2"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_DREPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: LPM_HINT STRING "LPM_REMAINDERPOSITIVE=TRUE"
// Retrieval info: CONSTANT: LPM_NREPRESENTATION STRING "SIGNED"
// Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "25"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_DIVIDE"
// Retrieval info: CONSTANT: LPM_WIDTHD NUMERIC "21"
// Retrieval info: CONSTANT: LPM_WIDTHN NUMERIC "33"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: denom 0 0 21 0 INPUT NODEFVAL "denom[20..0]"
// Retrieval info: USED_PORT: numer 0 0 33 0 INPUT NODEFVAL "numer[32..0]"
// Retrieval info: USED_PORT: quotient 0 0 33 0 OUTPUT NODEFVAL "quotient[32..0]"
// Retrieval info: USED_PORT: remain 0 0 21 0 OUTPUT NODEFVAL "remain[20..0]"
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @denom 0 0 21 0 denom 0 0 21 0
// Retrieval info: CONNECT: @numer 0 0 33 0 numer 0 0 33 0
// Retrieval info: CONNECT: quotient 0 0 33 0 @quotient 0 0 33 0
// Retrieval info: CONNECT: remain 0 0 21 0 @remain 0 0 21 0
// Retrieval info: GEN_FILE: TYPE_NORMAL div.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL div.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL div.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL div.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL div_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL div_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
